/********************
* Filename:		noc_router_tb.v
* Description:	Testbench for NOC Router Architecture with minimal functionality that contains the data path of 5 port(North, East, West, South, Local) 
                Input port FIFO buffer along with Control Path of LBDR and the arbiter. 
                Each Input port buffer has got LBDR routing module and the arbiter sends the grant coming from one of the LBDR 
                based on Round-Robin scheduling to the port decoder which asserts the respective read enable along with the 
                select lines to select the output port for the crossbar switch. 
                Active high control signals. Reset signal is active high synchronous reset
*
* $Revision: 36 $
* $Id: noc_router_tb.v 36 2016-02-20 16:43:26Z ranga $
* $Date: 2016-02-20 18:43:26 +0200 (Sat, 20 Feb 2016) $
* $Author: ranga $
*********************/
`timescale 1ns / 1ns
`include "../include/parameters.v"
`include "../include/state_defines.v"

module noc_router_tb;

/* 

 HEADER FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |         |         |        |       |   | 
   | 31 - 29  | 28 - 17 | 16 - 13 | 12 - 9 | 8 - 1 | 0 |
   |          |         |         |        |       |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE 			      (3 bits, one-hot encoded: Header=001)
 FLIT [28 : 17] = PACKET LENGTH         (12 bits, packet length in terms of # of flits = Header + Body (Payload) + Tail
 FLIT [16 : 13] = DESTINATION ADDRESS   (4 bits, addressing a 4x4 2D Mesh NoC at most)
 FLIT [12 : 9]  = SOURCE ADDRESS 	      (4 bits, addressing a 4x4 2D Mesh NoC at most)
 FLIT [8 : 1]   = PACKET ID        	    (ont-hot encoded counter, generated by NI, for ordering packets and flits in them)
 FLIT [0]       = PARITY BIT 			      (odd parity bit) 


 BODY (PAYLOAD) FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |                                    |   | 
   | 31 - 29  |                28 - 1              | 0 |
   |          |                                    |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE       (3 bits, one-hot encoded: Body (Payload)=010)
 FLIT [28 : 1]  = DATA (PAYLOAD)  (28 bits, actual data (payload) to be transmitted) 
 FLIT [0]       = PARITY BIT      (odd parity bit) 


 TAIL FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |                                    |   | 
   | 31 - 29  |                28 - 1              | 0 |
   |          |                                    |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE       (3 bits, one-hot encoded: Tail=100)
 FLIT [28 : 1]  = DATA (PAYLOAD)  (28 bits, actual data (Tail) to be transmitted)
 FLIT [0]       = PARITY BIT      (odd parity bit) 

*/
  
  // Declaring the port variables for DUT
  reg                      clk, rst;                                                         // rst is active low!
  reg [7:0]                Rxy;                                                              // Routing bits set during reset
  reg [3:0]                Cx;                                                               // Connectivity bits set during reset
  reg [`AXIS-1 : 0]   cur_addr;                                                         // currrent address of the router set during reset
  reg [`DATA_WIDTH-1 : 0]  Ldata_in, Ndata_in, Edata_in, Wdata_in, Sdata_in;                 // Incoming data from PREVIOUS router(NI)
  reg                      Lvalid_in, Nvalid_in, Evalid_in, Wvalid_in, Svalid_in;            // Incoming valid signal from PREVIOUS router(NI)
  reg                      Lready_in, Nready_in, Eready_in, Wready_in, Sready_in;            // Incoming ready signal from NEXT router(NI)
  
  wire [`DATA_WIDTH-1 : 0] Ldata_out, Ndata_out, Edata_out, Wdata_out, Sdata_out;            // Outgoing data to NEXT router(NI)
  wire                     Lready_out, Nready_out, Eready_out, Wready_out, Sready_out;       // Outgoing ready signal to PREVIOUS router(NI)
  wire                     Lvalid_out, Nvalid_out, Evalid_out, Wvalid_out, Svalid_out;       // Outgoing valid signal to NEXT router(NI)
  //wire                     Lparity_err, Nparity_err, Eparity_err, Wparity_err, Sparity_err;  // Parity error checker along with data_out
    
  // Instantiate NOC_ROUTER DUT
  noc_router DUT (clk, rst,
                  Rxy, Cx, cur_addr,
                  Ldata_in, Lvalid_in, Lready_out, Ldata_out, Lvalid_out, Lready_in,
                  Ndata_in, Nvalid_in, Nready_out, Ndata_out, Nvalid_out, Nready_in,
                  Edata_in, Evalid_in, Eready_out, Edata_out, Evalid_out, Eready_in,
                  Wdata_in, Wvalid_in, Wready_out, Wdata_out, Wvalid_out, Wready_in,
                  Sdata_in, Svalid_in, Sready_out, Sdata_out, Svalid_out, Sready_in/*,
                  Lparity_err, Nparity_err, Eparity_err, Wparity_err, Sparity_err*/
                );

  // Assertions 
  assert a0( .clk(clk), .valid(Nvalid_out), .data_out (Ndata_out));
  assert a1( .clk(clk), .valid(Evalid_out), .data_out (Edata_out));
  assert a2( .clk(clk), .valid(Wvalid_out), .data_out (Wdata_out));
  assert a3( .clk(clk), .valid(Svalid_out), .data_out (Sdata_out));
  assert a4( .clk(clk), .valid(Lvalid_out), .data_out (Ldata_out));
                  
  // Declaring the local variables
  reg [27 : 0]            data;               // 28 bits
  reg [2 : 0]             flit;
  reg                     parity = 1;
  reg [`DATA_WIDTH-1 : 0] tmp_data;
  
  `include "tb_tasks.v"             // to include task predefined after declaring the signals
  
  // Specify the CYCLE parameter
  parameter CYCLE = 10;
  
  // Generating Clock of period 10ns
  initial begin
    clk = 0;
    forever 
      #(CYCLE/2) clk = ~clk;
  end
  
  // Start the simulation
  initial begin : SIM
    integer i;
    
    // Reset & Initialize
    // reset(.Rxy_rst, .Cx_rst, .cur_addr_rst)
    // xpkt_gen(.p_length, .d_addr, .s_addr, .p_id);
/*  reset(8'b00111100, 4'b1110, 4'b0001); //--NODE1
    Npkt_gen(12'd10, 4'd8, 4'd1, 8'd1); // West
    #(CYCLE * 5);
    reset(8'b00111100, 4'b1111, 4'b1010); //--NODE10
    Epkt_gen(12'd5, 4'd14, 4'd5, 8'd2); // South
    #(CYCLE * 5); 
    reset(8'b00111100, 4'b1111, 4'b0101); //--NODE5
    Wpkt_gen(12'd20, 4'd5, 4'd14, 8'd3); // Local
    #(CYCLE * 5); 
    reset(8'b00111100, 4'b0101, 4'b1111); //--NODE15
    Spkt_gen(12'd3, 4'd3, 4'd12, 8'd4); // North
    #(CYCLE * 5); 
    reset(8'b00111100, 4'b1011, 4'b1000); //--NODE8
    Lpkt_gen(12'd7, 4'd11, 4'd8, 8'd5); // East
    #(CYCLE * 5); 
    reset(8'b00111100, 4'b1111, 4'b0101); //--NODE5
    fork
      Npkt_gen(12'd7, 4'd8, 4'd1, 8'd1); // West
      Epkt_gen(12'd12, 4'd14, 4'd5, 8'd2); // East
      Wpkt_gen(12'd4, 4'd5, 4'd14, 8'd3); // Local
      Spkt_gen(12'd20, 4'd3, 4'd12, 8'd4); // East
      Lpkt_gen(12'd8, 4'd11, 4'd8, 8'd5); // East
    join
*/

    reset(8'b00111100, 4'b1111, 4'b0101); //--NODE5
	// -----------------------------	 case: 1437
// -----------------------------	 case: 0

	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
#(4 * CYCLE);
// -----------------------------	 case: 1
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
#(4 * CYCLE);
// -----------------------------	 case: 2
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
#(4 * CYCLE);
// -----------------------------	 case: 3
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
#(4 * CYCLE);
// -----------------------------	 case: 4
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
#(4 * CYCLE);
// -----------------------------	 case: 5
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
#(4 * CYCLE);
// -----------------------------	 case: 6
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
#(4 * CYCLE);
// -----------------------------	 case: 7
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
#(4 * CYCLE);
// -----------------------------	 case: 8
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
#(4 * CYCLE);
// -----------------------------	 case: 9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
#(4 * CYCLE);
// -----------------------------	 case: 10
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
#(4 * CYCLE);
// -----------------------------	 case: 11
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
#(4 * CYCLE);
// -----------------------------	 case: 12
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
#(4 * CYCLE);
// -----------------------------	 case: 13
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd1); 	// E_W    6->0
#(4 * CYCLE);
// -----------------------------	 case: 14
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd1); 	// S_N    9->1
#(4 * CYCLE);
// -----------------------------	 case: 15
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd1); 	// N_S    1->9
#(4 * CYCLE);
// -----------------------------	 case: 16
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
join
#(4 * CYCLE);
// -----------------------------	 case: 17
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 18
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 19
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 20
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 21
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 22
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 23
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 24
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 25
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
join
#(4 * CYCLE);
// -----------------------------	 case: 26
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 27
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 28
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 29
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 30
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 31
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 32
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 33
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 34
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 35
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 36
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 37
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 38
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 39
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 40
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 41
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 42
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 43
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 44
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 45
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 46
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 47
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 48
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 49
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 50
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 51
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 52
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 53
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 54
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 55
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 56
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 57
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 58
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 59
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 60
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 61
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 62
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 63
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 64
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 65
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 66
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 67
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 68
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 69
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 70
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 71
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 72
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 73
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 74
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 75
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 76
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 77
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 78
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 79
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 80
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 81
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 82
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 83
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 84
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 85
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 86
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 87
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 88
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 89
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 90
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 91
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 92
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 93
fork
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd1); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 94
fork
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd1); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 95
fork
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd1); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 96
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 97
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 98
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 99
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 100
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 101
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 102
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 103
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 104
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 105
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 106
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 107
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 108
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 109
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 110
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 111
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 112
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 113
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 114
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 115
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 116
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 117
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 118
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 119
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 120
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 121
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 122
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 123
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 124
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 125
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 126
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 127
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 128
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 129
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 130
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 131
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 132
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 133
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 134
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 135
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 136
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 137
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 138
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 139
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 140
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 141
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 142
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 143
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 144
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 145
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 146
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 147
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 148
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 149
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 150
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 151
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 152
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 153
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 154
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 155
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 156
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 157
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 158
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 159
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 160
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 161
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 162
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 163
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 164
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 165
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 166
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 167
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 168
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 169
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 170
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 171
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 172
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 173
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 174
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 175
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 176
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 177
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 178
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 179
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 180
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 181
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 182
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 183
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 184
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 185
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 186
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 187
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 188
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 189
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 190
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 191
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 192
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 193
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 194
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 195
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 196
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 197
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 198
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 199
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 200
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 201
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 202
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 203
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 204
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 205
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 206
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 207
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 208
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 209
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 210
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 211
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 212
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 213
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 214
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 215
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 216
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 217
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 218
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 219
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 220
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 221
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 222
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 223
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 224
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 225
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 226
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 227
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 228
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 229
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 230
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 231
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 232
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 233
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 234
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 235
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 236
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 237
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 238
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 239
fork
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd1); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 240
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 241
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 242
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 243
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 244
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 245
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 246
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 247
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 248
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 249
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 250
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 251
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 252
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 253
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 254
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 255
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 256
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 257
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 258
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 259
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 260
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 261
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 262
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 263
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 264
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 265
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 266
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 267
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 268
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 269
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 270
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 271
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 272
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 273
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 274
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 275
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 276
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 277
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 278
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 279
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 280
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 281
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 282
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 283
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 284
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 285
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 286
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 287
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 288
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 289
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 290
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 291
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 292
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 293
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 294
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 295
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 296
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 297
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 298
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 299
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 300
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 301
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 302
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 303
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 304
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 305
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 306
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 307
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 308
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 309
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 310
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 311
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 312
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 313
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 314
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 315
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 316
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 317
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 318
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 319
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 320
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 321
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 322
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 323
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 324
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 325
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 326
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 327
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 328
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 329
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
join
#(4 * CYCLE);
// -----------------------------	 case: 330
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
join
#(4 * CYCLE);
// -----------------------------	 case: 331
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 332
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 333
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 334
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 335
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 336
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 337
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 338
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 339
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 340
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 341
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
join
#(4 * CYCLE);
// -----------------------------	 case: 342
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 343
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 344
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 345
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 346
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 347
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 348
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 349
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 350
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 351
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 352
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
join
#(4 * CYCLE);
// -----------------------------	 case: 353
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 354
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 355
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 356
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 357
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 358
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 359
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 360
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 361
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 362
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 363
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 364
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 365
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 366
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 367
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 368
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 369
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 370
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 371
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 372
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 373
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 374
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 375
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 376
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 377
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 378
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 379
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 380
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 381
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 382
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 383
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 384
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 385
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 386
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 387
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 388
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 389
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 390
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 391
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 392
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 393
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 394
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 395
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 396
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 397
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 398
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 399
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 400
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 401
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 402
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 403
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 404
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 405
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 406
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 407
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 408
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 409
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 410
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 411
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 412
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 413
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 414
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 415
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 416
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 417
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 418
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 419
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 420
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 421
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 422
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 423
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 424
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 425
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 426
fork
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd1); 	// E_W    6->0
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 427
fork
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd1); 	// E_W    6->0
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 428
fork
	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd1); 	// S_N    9->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd2); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 429
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 430
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 431
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 432
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 433
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 434
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 435
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 436
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 437
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 438
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 439
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 440
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 441
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 442
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 443
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 444
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 445
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 446
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 447
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 448
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 449
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 450
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 451
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 452
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 453
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 454
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 455
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 456
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 457
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 458
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 459
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 460
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 461
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 462
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 463
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 464
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 465
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 466
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 467
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 468
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 469
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 470
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 471
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 472
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 473
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 474
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 475
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 476
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 477
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 478
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 479
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 480
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 481
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 482
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 483
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 484
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 485
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 486
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 487
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 488
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 489
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 490
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 491
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 492
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 493
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 494
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 495
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 496
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 497
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 498
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 499
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 500
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 501
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 502
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 503
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 504
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 505
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 506
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 507
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 508
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 509
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 510
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 511
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 512
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 513
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 514
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 515
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 516
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 517
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 518
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 519
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 520
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 521
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 522
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 523
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 524
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 525
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
join
#(4 * CYCLE);
// -----------------------------	 case: 526
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
join
#(4 * CYCLE);
// -----------------------------	 case: 527
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
join
#(4 * CYCLE);
// -----------------------------	 case: 528
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
join
#(4 * CYCLE);
// -----------------------------	 case: 529
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 530
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 531
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 532
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 533
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 534
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 535
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 536
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 537
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 538
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 539
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 540
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 541
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 542
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 543
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 544
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 545
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 546
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 547
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 548
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 549
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 550
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 551
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 552
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 553
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 554
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 555
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 556
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 557
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 558
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 559
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 560
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 561
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 562
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 563
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 564
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 565
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 566
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 567
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 568
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 569
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 570
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 571
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 572
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 573
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 574
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 575
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 576
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 577
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 578
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 579
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 580
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 581
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 582
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 583
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 584
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 585
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 586
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 587
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
join
#(4 * CYCLE);
// -----------------------------	 case: 588
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 589
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 590
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 591
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 592
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 593
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 594
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 595
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 596
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 597
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 598
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 599
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 600
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 601
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 602
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 603
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 604
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 605
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 606
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 607
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 608
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 609
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 610
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 611
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 612
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 613
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 614
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 615
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 616
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 617
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 618
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 619
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 620
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 621
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 622
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 623
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 624
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 625
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 626
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 627
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 628
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 629
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 630
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 631
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 632
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 633
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 634
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 635
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 636
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 637
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 638
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 639
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 640
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 641
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 642
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 643
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 644
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 645
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 646
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 647
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 648
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 649
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 650
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 651
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 652
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 653
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 654
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 655
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 656
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 657
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 658
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 659
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 660
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 661
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 662
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 663
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 664
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 665
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 666
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 667
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 668
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 669
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 670
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 671
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 672
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 673
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 674
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 675
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 676
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 677
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 678
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 679
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 680
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 681
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 682
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 683
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 684
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 685
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 686
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 687
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 688
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 689
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 690
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 691
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 692
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 693
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 694
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 695
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 696
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 697
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 698
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 699
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 700
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 701
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 702
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 703
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 704
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 705
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 706
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 707
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 708
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 709
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 710
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 711
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 712
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 713
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 714
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 715
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 716
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 717
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 718
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 719
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 720
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 721
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 722
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 723
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 724
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 725
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 726
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 727
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 728
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 729
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 730
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 731
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 732
fork
	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd1); 	// E_W    6->0
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd2); 	// S_N    9->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd3); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 733
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 734
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 735
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 736
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 737
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 738
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 739
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 740
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 741
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 742
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 743
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 744
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 745
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 746
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 747
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 748
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 749
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 750
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 751
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 752
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 753
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 754
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 755
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 756
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 757
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 758
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 759
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 760
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 761
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 762
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 763
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 764
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 765
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 766
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 767
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 768
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 769
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 770
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 771
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 772
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 773
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 774
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 775
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 776
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 777
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 778
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 779
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 780
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 781
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 782
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 783
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 784
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 785
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 786
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 787
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 788
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 789
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 790
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 791
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 792
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 793
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 794
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 795
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 796
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 797
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 798
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 799
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 800
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 801
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 802
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 803
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 804
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 805
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 806
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 807
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 808
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 809
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 810
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 811
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 812
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 813
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 814
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 815
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 816
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 817
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 818
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 819
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 820
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 821
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 822
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 823
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 824
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 825
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 826
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 827
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 828
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 829
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 830
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 831
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 832
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 833
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 834
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 835
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 836
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 837
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 838
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 839
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 840
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 841
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 842
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 843
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 844
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 845
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 846
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 847
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 848
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 849
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 850
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 851
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 852
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 853
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 854
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 855
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 856
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 857
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 858
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 859
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 860
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 861
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 862
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 863
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 864
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 865
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 866
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 867
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 868
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 869
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 870
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 871
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 872
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 873
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 874
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 875
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 876
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 877
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 878
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 879
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 880
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 881
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 882
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 883
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 884
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 885
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 886
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 887
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 888
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 889
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 890
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 891
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 892
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 893
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 894
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 895
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 896
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 897
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 898
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 899
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 900
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 901
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 902
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 903
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 904
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 905
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 906
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 907
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 908
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 909
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 910
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 911
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 912
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 913
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 914
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 915
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 916
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 917
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 918
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 919
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 920
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 921
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 922
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 923
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 924
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 925
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 926
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 927
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 928
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 929
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 930
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 931
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 932
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 933
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 934
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 935
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 936
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 937
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 938
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 939
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 940
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 941
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 942
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 943
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 944
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 945
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 946
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 947
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 948
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 949
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 950
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 951
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 952
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 953
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 954
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 955
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 956
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 957
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 958
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 959
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 960
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 961
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 962
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 963
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 964
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 965
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 966
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 967
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 968
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 969
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 970
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 971
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 972
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 973
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 974
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 975
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 976
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 977
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 978
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 979
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 980
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 981
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 982
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 983
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 984
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 985
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 986
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 987
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 988
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 989
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 990
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 991
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 992
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 993
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 994
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 995
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 996
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 997
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 998
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 999
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1000
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1001
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1002
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1003
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1004
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1005
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1006
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1007
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1008
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1009
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1010
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1011
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1012
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1013
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1014
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1015
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1016
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1017
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1018
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1019
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1020
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1021
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1022
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1023
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1024
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1025
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1026
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1027
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1028
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1029
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1030
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1031
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1032
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1033
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1034
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1035
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1036
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1037
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1038
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1039
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1040
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1041
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1042
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1043
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1044
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1045
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1046
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1047
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1048
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1049
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1050
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1051
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1052
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1053
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1054
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1055
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1056
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1057
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1058
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1059
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1060
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1061
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1062
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1063
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1064
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1065
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1066
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1067
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1068
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1069
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1070
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1071
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1072
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1073
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1074
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1075
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1076
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1077
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1078
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1079
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1080
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1081
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1082
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1083
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1084
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1085
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1086
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1087
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1088
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1089
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1090
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1091
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1092
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1093
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1094
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1095
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1096
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1097
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1098
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1099
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1100
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1101
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1102
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1103
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1104
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1105
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1106
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1107
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1108
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1109
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1110
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1111
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1112
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1113
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1114
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1115
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1116
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1117
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1118
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1119
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1120
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1121
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1122
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1123
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1124
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1125
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1126
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1127
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1128
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1129
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1130
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1131
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1132
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1133
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1134
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1135
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1136
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1137
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1138
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1139
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1140
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1141
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1142
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1143
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1144
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1145
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1146
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1147
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1148
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1149
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1150
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1151
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1152
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1153
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1154
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1155
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1156
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1157
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1158
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1159
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1160
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1161
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1162
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1163
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1164
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1165
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1166
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1167
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1168
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1169
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1170
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1171
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1172
fork
	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd1); 	// E2L    6->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1173
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1174
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1175
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1176
fork
	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd1); 	// N2L    1->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1177
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1178
fork
	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd1); 	// W2L    4->5
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1179
fork
	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd1); 	// S2L    9->5
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1180
fork
	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd1); 	// W_E    4->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd2); 	// E_W    6->0
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd3); 	// S_N    9->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd4); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1181
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1182
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1183
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1184
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1185
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1186
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1187
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1188
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1189
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1190
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1191
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1192
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1193
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1194
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1195
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1196
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd2); 	// W2N    4->1
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1197
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1198
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1199
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1200
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1201
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1202
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1203
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1204
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1205
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1206
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1207
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1208
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1209
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1210
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1211
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1212
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1213
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1214
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1215
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1216
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1217
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1218
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1219
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1220
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1221
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1222
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1223
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1224
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1225
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1226
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1227
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1228
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1229
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1230
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1231
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1232
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1233
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1234
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1235
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1236
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1237
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1238
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1239
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1240
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1241
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1242
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1243
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1244
fork
	Epkt_gen(12'd12, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1245
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1246
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1247
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1248
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1249
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1250
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1251
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1252
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1253
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1254
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1255
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1256
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1257
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1258
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1259
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1260
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd2); 	// E2S    6->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1261
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1262
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1263
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1264
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1265
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1266
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1267
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1268
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1269
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1270
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1271
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1272
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1273
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1274
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1275
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1276
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1277
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1278
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1279
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1280
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1281
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1282
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1283
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1284
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1285
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1286
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1287
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1288
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1289
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1290
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1291
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1292
fork
	Wpkt_gen(12'd12, 4'd1, 4'd4, 8'd1); 	// W2N    4->1
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1293
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1294
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1295
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1296
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd3); 	// L2E    5->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1297
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1298
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1299
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1300
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd3); 	// L2N    5->1
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1301
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1302
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1303
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1304
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1305
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1306
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1307
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1308
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd2); 	// W2S    4->9
	#(2*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd3); 	// L2W    5->4
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1309
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1310
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1311
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1312
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1313
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1314
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1315
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1316
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1317
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1318
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1319
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1320
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1321
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1322
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1323
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1324
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1325
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1326
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1327
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1328
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1329
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1330
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1331
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1332
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1333
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1334
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1335
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1336
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1337
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1338
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1339
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1340
fork
	Epkt_gen(12'd12, 4'd9, 4'd6, 8'd1); 	// E2S    6->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1341
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1342
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1343
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1344
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1345
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1346
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1347
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1348
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd2); 	// L2E    5->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1349
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1350
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1351
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1352
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1353
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1354
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1355
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1356
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1357
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1358
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1359
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1360
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1361
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1362
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1363
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1364
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd2); 	// L2S    5->9
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1365
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1366
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd4); 	// N2L    1->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1367
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1368
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd3); 	// E2L    6->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1369
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1370
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1371
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1372
fork
	Wpkt_gen(12'd12, 4'd9, 4'd4, 8'd1); 	// W2S    4->9
	#(1*CYCLE)	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd2); 	// L2W    5->4
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1373
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1374
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1375
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1376
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1377
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1378
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1379
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1380
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1381
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1382
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1383
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1384
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1385
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1386
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1387
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1388
fork
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1389
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1390
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1391
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1392
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1393
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1394
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1395
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1396
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1397
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1398
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1399
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1400
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1401
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1402
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1403
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1404
fork
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd1); 	// L2N    5->1
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1405
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1406
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1407
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1408
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1409
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1410
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1411
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1412
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1413
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1414
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1415
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1416
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1417
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1418
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1419
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1420
fork
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd1); 	// L2S    5->9
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1421
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd5); 	// S2L    9->5
join
#(4 * CYCLE);
// -----------------------------	 case: 1422
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd4); 	// W2L    4->5
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1423
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd5); 	// W_E    4->6
join
#(4 * CYCLE);
// -----------------------------	 case: 1424
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd3); 	// N2L    1->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1425
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1426
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1427
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1428
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Epkt_gen(12'd12, 4'd5, 4'd6, 8'd2); 	// E2L    6->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1429
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd4); 	// S2L    9->5
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1430
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd3); 	// W2L    4->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1431
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd4); 	// W_E    4->6
	#(4*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd5); 	// E_W    6->0
join
#(4 * CYCLE);
// -----------------------------	 case: 1432
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Npkt_gen(12'd12, 4'd5, 4'd1, 8'd2); 	// N2L    1->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd5); 	// S_N    9->1
join
#(4 * CYCLE);
// -----------------------------	 case: 1433
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd3); 	// S2L    9->5
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1434
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd5, 4'd4, 8'd2); 	// W2L    4->5
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1435
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Spkt_gen(12'd12, 4'd5, 4'd9, 8'd2); 	// S2L    9->5
	#(2*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd3); 	// W_E    4->6
	#(3*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd4); 	// E_W    6->0
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1436
fork
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd1); 	// L2W    5->4
	#(1*CYCLE)	Wpkt_gen(12'd12, 4'd6, 4'd4, 8'd2); 	// W_E    4->6
	#(2*CYCLE)	Epkt_gen(12'd12, 4'd0, 4'd6, 8'd3); 	// E_W    6->0
	#(3*CYCLE)	Spkt_gen(12'd12, 4'd1, 4'd9, 8'd4); 	// S_N    9->1
	#(4*CYCLE)	Npkt_gen(12'd12, 4'd9, 4'd1, 8'd5); 	// N_S    1->9
join
#(4 * CYCLE);
// -----------------------------	 case: 1437
	Lpkt_gen(12'd12, 4'd6, 4'd5, 8'd1); 	// L2E    5->6
	Lpkt_gen(12'd12, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	Lpkt_gen(12'd12, 4'd9, 4'd5, 8'd3); 	// L2S    5->9
	Lpkt_gen(12'd12, 4'd4, 4'd5, 8'd4); 	// L2W    5->4


#(4 * CYCLE);

	fork
	Lpkt_gen(12'd5, 4'd1, 4'd5, 8'd2); 	// L2N    5->1
	#(3*CYCLE) Epkt_gen(12'd5, 4'd1, 4'd6, 8'd1); 	// E2N    6->1
	join
    #(CYCLE * 25);
    $stop;
  end

  initial begin
    $monitor("TIME:%0t *********STATUS:: Ldata_out:%0h, Ndata_out:%0h, Edata_out:%0h, Wdata_out:%0h, Sdata_out:%0h, Lready_out:%0b, Nready_out:%0b, Eready_out:%0b, Wready_out:%0b, Sready_out:%0b,  Lvalid_out:%0b, Nvalid_out:%0b, Evalid_out:%0b, Wvalid_out:%0b, Svalid_out:%0b", $time, Ldata_out, Ndata_out, Edata_out, Wdata_out, Sdata_out, Lready_out, Nready_out, Eready_out, Wready_out, Sready_out, Lvalid_out, Nvalid_out, Evalid_out, Wvalid_out, Svalid_out);
  end

endmodule

module assert(input clk, input valid, input [31 : 0] data_out);
 
//    integer f;
integer packet_started = 0; // boolean value

    always @(posedge clk)
    begin
	if ( packet_started == 1 && (data_out[(`DATA_WIDTH-1) : (`DATA_WIDTH-3)] == 0'b001)) // HEADER flit
	    begin
	       $display("TIME: %0t Error!\n", $time);
	       $stop;
	end
	if (valid == 1) // ?? This means when the packet is sent until the end
        begin
	    
	    if ( data_out[(`DATA_WIDTH-1) : (`DATA_WIDTH-3)] == 0'b001) // HEADER flit
	    begin
	       packet_started = 1;
	    end
	    if ( data_out[(`DATA_WIDTH-1) : (`DATA_WIDTH-3)] == 0'b100) // TAIL flit
	    begin
	       packet_started = 0;
	    end
	end
    end

    always @(data_out)
    begin
        if (valid == 1) // ?? This means when the packet is sent until the end
        begin
	//    f = $fopen("output.txt","a");
//	    $fdisplay(f,"TIME: %0t FLIT_TYPE: %0b DST_ADDR: %0b \n", $time, data_out[(`DATA_WIDTH-19) +: 2]);
            $display("Received: TIME: %0t FLIT_TYPE: %0b DST_ADDR: %0b \n", $time,  data_out[(`DATA_WIDTH-1) : (`DATA_WIDTH-3)], data_out[28 : 25]);
//	    $fclose(f);
	   
     
	    
        end
    end
endmodule

