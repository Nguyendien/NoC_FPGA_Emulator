/********************
* Filename:		noc_router_tb.v
* Description:	Testbench for NOC Router Architecture with minimal functionality that contains the data path of 5 port(North, East, West, South, Local) 
                Input port FIFO buffer along with Control Path of LBDR and the arbiter. 
                Each Input port buffer has got LBDR routing module and the arbiter sends the grant coming from one of the LBDR 
                based on Round-Robin scheduling to the port decoder which asserts the respective read enable along with the 
                select lines to select the output port for the crossbar switch. 
                Active high control signals. Reset signal is active high synchronous reset
*
* $Revision: 36 $
* $Id: noc_router_tb.v 36 2016-02-20 16:43:26Z ranga $
* $Date: 2016-02-20 18:43:26 +0200 (Sat, 20 Feb 2016) $
* $Author: ranga $
*********************/
`include "../include/parameters.v"
`include "../include/state_defines.v"

module noc_router_tb;

/* 

 HEADER FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |         |         |        |       |   | 
   | 31 - 29  | 28 - 17 | 16 - 13 | 12 - 9 | 8 - 1 | 0 |
   |          |         |         |        |       |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE 			      (3 bits, one-hot encoded: Header=001)
 FLIT [28 : 17] = PACKET LENGTH         (12 bits, packet length in terms of # of flits = Header + Body (Payload) + Tail
 FLIT [16 : 13] = DESTINATION ADDRESS   (4 bits, addressing a 4x4 2D Mesh NoC at most)
 FLIT [12 : 9]  = SOURCE ADDRESS 	      (4 bits, addressing a 4x4 2D Mesh NoC at most)
 FLIT [8 : 1]   = PACKET ID        	    (ont-hot encoded counter, generated by NI, for ordering packets and flits in them)
 FLIT [0]       = PARITY BIT 			      (odd parity bit) 


 BODY (PAYLOAD) FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |                                    |   | 
   | 31 - 29  |                28 - 1              | 0 |
   |          |                                    |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE       (3 bits, one-hot encoded: Body (Payload)=010)
 FLIT [28 : 1]  = DATA (PAYLOAD)  (28 bits, actual data (payload) to be transmitted) 
 FLIT [0]       = PARITY BIT      (odd parity bit) 


 TAIL FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |                                    |   | 
   | 31 - 29  |                28 - 1              | 0 |
   |          |                                    |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE       (3 bits, one-hot encoded: Tail=100)
 FLIT [28 : 1]  = DATA (PAYLOAD)  (28 bits, actual data (Tail) to be transmitted)
 FLIT [0]       = PARITY BIT      (odd parity bit) 

*/
  
  // Declaring the port variables for DUT
  reg                      clk, rst;
  reg [7:0]                Rxy;                                                              // Routing bits set during reset
  reg [3:0]                Cx;                                                               // Connectivity bits set during reset
  reg [`AXIS-1 : 0]   cur_addr;                                                         // currrent address of the router set during reset
  reg [`DATA_WIDTH-1 : 0]  Ldata_in, Ndata_in, Edata_in, Wdata_in, Sdata_in;                 // Incoming data from PREVIOUS router(NI)
  reg                      Lvalid_in, Nvalid_in, Evalid_in, Wvalid_in, Svalid_in;            // Incoming valid signal from PREVIOUS router(NI)
  reg                      Lready_in, Nready_in, Eready_in, Wready_in, Sready_in;            // Incoming ready signal from NEXT router(NI)
  
  wire [`DATA_WIDTH-1 : 0] Ldata_out, Ndata_out, Edata_out, Wdata_out, Sdata_out;            // Outgoing data to NEXT router(NI)
  wire                     Lready_out, Nready_out, Eready_out, Wready_out, Sready_out;       // Outgoing ready signal to PREVIOUS router(NI)
  wire                     Lvalid_out, Nvalid_out, Evalid_out, Wvalid_out, Svalid_out;       // Outgoing valid signal to NEXT router(NI)
  //wire                     Lparity_err, Nparity_err, Eparity_err, Wparity_err, Sparity_err;  // Parity error checker along with data_out
    
  // Instantiate NOC_ROUTER DUT
  noc_router DUT (clk, rst,
                  Rxy, Cx, cur_addr,
                  Ldata_in, Lvalid_in, Lready_out, Ldata_out, Lvalid_out, Lready_in,
                  Ndata_in, Nvalid_in, Nready_out, Ndata_out, Nvalid_out, Nready_in,
                  Edata_in, Evalid_in, Eready_out, Edata_out, Evalid_out, Eready_in,
                  Wdata_in, Wvalid_in, Wready_out, Wdata_out, Wvalid_out, Wready_in,
                  Sdata_in, Svalid_in, Sready_out, Sdata_out, Svalid_out, Sready_in/*,
                  Lparity_err, Nparity_err, Eparity_err, Wparity_err, Sparity_err*/
                );
                  
  // Declaring the local variables
  reg [27 : 0]            data;               // 28 bits
  reg [2 : 0]             flit;
  reg                     parity = 1;
  reg [`DATA_WIDTH-1 : 0] tmp_data;
  
  `include "tb_tasks.v"             // to include task predefined after declaring the signals
  
  // Specify the CYCLE parameter
  parameter CYCLE = 10;
  
  // Generating Clock of period 10ns
  initial begin
    clk = 0;
    forever 
      #(CYCLE/2) clk = ~clk;
  end
  
  // Start the simulation
  initial begin : SIM
    integer i;
    
    // Reset & Initialize
    // reset(.Rxy_rst, .Cx_rst, .cur_addr_rst)
    // xpkt_gen(.p_length, .d_addr, .s_addr, .p_id);
    reset(8'b00111100, 4'b1110, 4'b0001); //--NODE1
    Npkt_gen(12'd10, 4'd8, 4'd1, 8'd1); // West
    #(CYCLE * 5);
    reset(8'b00111100, 4'b1111, 4'b1010); //--NODE10
    Epkt_gen(12'd5, 4'd14, 4'd5, 8'd2); // South
    #(CYCLE * 5); 
    reset(8'b00111100, 4'b1111, 4'b0101); //--NODE5
    Wpkt_gen(12'd20, 4'd5, 4'd14, 8'd3); // Local
    #(CYCLE * 5); 
    reset(8'b00111100, 4'b0101, 4'b1111); //--NODE15
    Spkt_gen(12'd3, 4'd3, 4'd12, 8'd4); // North
    #(CYCLE * 5); 
    reset(8'b00111100, 4'b1011, 4'b1000); //--NODE8
    Lpkt_gen(12'd7, 4'd11, 4'd8, 8'd5); // East
    #(CYCLE * 5); 
    reset(8'b00111100, 4'b1111, 4'b0101); //--NODE5
    fork
      Npkt_gen(12'd7, 4'd8, 4'd1, 8'd1); // West
      Epkt_gen(12'd12, 4'd14, 4'd5, 8'd2); // East
      Wpkt_gen(12'd4, 4'd5, 4'd14, 8'd3); // Local
      Spkt_gen(12'd20, 4'd3, 4'd12, 8'd4); // East
      Lpkt_gen(12'd8, 4'd11, 4'd8, 8'd5); // East
    join
    #(CYCLE * 25);
    $finish;
  end

  initial begin
    $monitor("TIME:%0t *********STATUS:: Ldata_out:%0h, Ndata_out:%0h, Edata_out:%0h, Wdata_out:%0h, Sdata_out:%0h, Lready_out:%0b, Nready_out:%0b, Eready_out:%0b, Wready_out:%0b, Sready_out:%0b,  Lvalid_out:%0b, Nvalid_out:%0b, Evalid_out:%0b, Wvalid_out:%0b, Svalid_out:%0b", $time, Ldata_out, Ndata_out, Edata_out, Wdata_out, Sdata_out, Lready_out, Nready_out, Eready_out, Wready_out, Sready_out, Lvalid_out, Nvalid_out, Evalid_out, Wvalid_out, Svalid_out);
  end

endmodule