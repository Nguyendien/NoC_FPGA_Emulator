/********************
* Filename:		noc_network_tb.v
* Description:	Testbench for NOC Network Architecture with minimal functionality that contains the data path of 5 port(North, East, West, South, Local) 
                2x2 Mesh Network
*
* $Revision: 39 $
* $Id: noc_network_tb.v 39 2016-02-20 19:11:39Z ranga $
* $Date: 2016-02-20 21:11:39 +0200 (Sat, 20 Feb 2016) $
* $Author: ranga $
*********************/
`include "../include/parameters.v"
`include "../include/state_defines.v"

module noc_network_tb;

/* 

 HEADER FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |         |         |        |       |   | 
   | 31 - 29  | 28 - 17 | 16 - 13 | 12 - 9 | 8 - 1 | 0 |
   |          |         |         |        |       |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE 			      (3 bits, one-hot encoded: Header=001)
 FLIT [28 : 17] = PACKET LENGTH         (12 bits, packet length in terms of # of flits = Header + Body (Payload) + Tail
 FLIT [16 : 13] = DESTINATION ADDRESS   (4 bits, addressing a 4x4 2D Mesh NoC at most)
 FLIT [12 : 9]  = SOURCE ADDRESS 	      (4 bits, addressing a 4x4 2D Mesh NoC at most)
 FLIT [8 : 1]   = PACKET ID        	    (ont-hot encoded counter, generated by NI, for ordering packets and flits in them)
 FLIT [0]       = PARITY BIT 			      (odd parity bit) 


 BODY (PAYLOAD) FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |                                    |   | 
   | 31 - 29  |                28 - 1              | 0 |
   |          |                                    |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE       (3 bits, one-hot encoded: Body (Payload)=010)
 FLIT [28 : 1]  = DATA (PAYLOAD)  (28 bits, actual data (payload) to be transmitted) 
 FLIT [0]       = PARITY BIT      (odd parity bit) 


 TAIL FLIT DESCRIPTION (32 bits - compatible with LEON3)
    ---------------------------------------------------
   |          |                                    |   | 
   | 31 - 29  |                28 - 1              | 0 |
   |          |                                    |   |
    ---------------------------------------------------

 FLIT [31 : 29] = FLIT TYPE       (3 bits, one-hot encoded: Tail=100)
 FLIT [28 : 1]  = DATA (PAYLOAD)  (28 bits, actual data (Tail) to be transmitted)
 FLIT [0]       = PARITY BIT      (odd parity bit) 

*/
  
  // Declaring the port variables for DUT
  reg                      clk, rst;
  reg [7:0]                Rxy[`NODES-1 : 0];                                                              // Routing bits set during reset
  reg [3:0]                Cx[`NODES-1 : 0];                                                               // Connectivity bits set during reset
  reg [`AXIS-1 : 0]   cur_addr[`NODES-1 : 0];                                                         // currrent address of the router set during reset
  reg [`DATA_WIDTH-1 : 0]  Ldata_in[`NODES-1 : 0], Ndata_in[`NODES-1 : 0], Edata_in[`NODES-1 : 0], Wdata_in[`NODES-1 : 0], Sdata_in[`NODES-1 : 0];                 // Incoming data from PREVIOUS router(NI)
  reg                      Lvalid_in[`NODES-1 : 0], Nvalid_in[`NODES-1 : 0], Evalid_in[`NODES-1 : 0], Wvalid_in[`NODES-1 : 0], Svalid_in[`NODES-1 : 0];            // Incoming valid signal from PREVIOUS router(NI)
  reg                      Lready_in[`NODES-1 : 0], Nready_in[`NODES-1 : 0], Eready_in[`NODES-1 : 0], Wready_in[`NODES-1 : 0], Sready_in[`NODES-1 : 0];            // Incoming ready signal from NEXT router(NI)
  
  wire [`DATA_WIDTH-1 : 0] Ldata_out[`NODES-1 : 0], Ndata_out[`NODES-1 : 0], Edata_out[`NODES-1 : 0], Wdata_out[`NODES-1 : 0], Sdata_out[`NODES-1 : 0];            // Outgoing data to NEXT router(NI)
  wire                     Lready_out[`NODES-1 : 0], Nready_out[`NODES-1 : 0], Eready_out[`NODES-1 : 0], Wready_out[`NODES-1 : 0], Sready_out[`NODES-1 : 0];       // Outgoing ready signal to PREVIOUS router(NI)
  wire                     Lvalid_out[`NODES-1 : 0], Nvalid_out[`NODES-1 : 0], Evalid_out[`NODES-1 : 0], Wvalid_out[`NODES-1 : 0], Svalid_out[`NODES-1 : 0];       // Outgoing valid signal to NEXT router(NI)
      
  // Instantiate NOC_ROUTER based on number of nodes 
  generate
    genvar i, j;
      for(i = 0; i < `NODES; i = i+1) begin
      	  for(i = 0; j < `NODES; j = j+1) begin
      	  
			   if (i == 0 && j == 0)
  			   		noc_router_NW ROUTER (clk, rst,
                            Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            );
                            
		       else if (i ==  `NODES - 1 && j == 0)
		       		noc_router_NE ROUTER (clk, rst,
                            Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            );
                            
		       else if (i == 0 && j == `NODES - 1)
		       	    noc_router_SW ROUTER (clk, rst,
                            Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            );
                            
		       else if (i == `NODES - 1 && j == `NODES - 1)
		            noc_router_SE ROUTER (clk, rst,
                            Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            );
                            
		       else if (i == 0)
		       		noc_router_N ROUTER (clk, rst,
                            Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            );
		       		
		       else if (i == `NODES - 1)
		       		noc_router_S ROUTER (clk, rst,
                            Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            );
                            
		       else if (j == 0)
		    		noc_router_W ROUTER (clk, rst,
                            Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            );
                            
		       else if (j == `NODES - 1)
		       		noc_router_E ROUTER (clk, rst,
                            Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            );
                            
		       else
		       
		       		noc_router_FULL ROUTER (Rxy[j * `NODES + i], Cx[j * `NODES + i], cur_addr[j * `NODES + i],
                            Ldata_in[j * `NODES + i], Lvalid_in[j * `NODES + i], Lready_out[j * `NODES + i], Ldata_out[j * `NODES + i], Lvalid_out[j * `NODES + i], Lready_in[j * `NODES + i],
                            Ndata_in[j * `NODES + i], Nvalid_in[j * `NODES + i], Nready_out[j * `NODES + i], Ndata_out[j * `NODES + i], Nvalid_out[j * `NODES + i], Nready_in[j * `NODES + i],
                            Edata_in[j * `NODES + i], Evalid_in[j * `NODES + i], Eready_out[j * `NODES + i], Edata_out[j * `NODES + i], Evalid_out[j * `NODES + i], Eready_in[j * `NODES + i],
                            Wdata_in[j * `NODES + i], Wvalid_in[j * `NODES + i], Wready_out[j * `NODES + i], Wdata_out[j * `NODES + i], Wvalid_out[j * `NODES + i], Wready_in[j * `NODES + i],
                            Sdata_in[j * `NODES + i], Svalid_in[j * `NODES + i], Sready_out[j * `NODES + i], Sdata_out[j * `NODES + i], Svalid_out[j * `NODES + i], Sready_in[j * `NODES + i]
                            ); 
		       		   		 	 
  			   end

      	 end
      end
  endgenerate
  
  // output connectivity
  always @(*) begin
  	integer i,j; 
  	      for(i = 0; i < `NODES; i = i+1) begin
      	  	for(i = 0; j < `NODES; j = j+1) begin
				
				if (i == 0 && j == 0)  // Router NW
				begin
					Wdata_in[j * `NODES + i + 1]  = Edata_out[j * `NODES + i];
    				Wvalid_in[j * `NODES + i + 1] = Evalid_out[0];
    				Eready_in[j * `NODES + i] = Wready_out[j * `NODES + i + 1];
    				Ndata_in[(j + 1) * `NODES + i]  = Sdata_out[j * `NODES + i];
    				Nvalid_in[(j + 1) * `NODES + i] = Svalid_out[j * `NODES + i];
    				Sready_in[j * `NODES + i] = Nready_out[(j + 1) * `NODES + i];
				end 
					
				else if (i == `NODES - 1 && j == 0)  // Router NE
				begin
					Edata_in[j * `NODES + i - 1]  = Wdata_out[j * `NODES + i];
    				Evalid_in[j * `NODES + i - 1] = Wvalid_out[j * `NODES + i];
				    Wready_in[j * `NODES + i] = Eready_out[j * `NODES + i - 1];
  		  		    Ndata_in[(j + 1) * `NODES + i]  = Sdata_out[j * `NODES + i];
  				    Nvalid_in[(j + 1) * `NODES + i] = Svalid_out[j * `NODES + i];
   				    Sready_in[j * `NODES + i] = Nready_out[(j + 1) * `NODES + i];
				end
				
				else if (i == `NODES - 1 && j == 0)  // Router SW
				begin
    				Wdata_in[3]  = Edata_out[2];
    				Wvalid_in[3] = Evalid_out[2];
    				Eready_in[2] = Wready_out[3];
    				Sdata_in[0]  = Ndata_out[2];
    				Svalid_in[0] = Nvalid_out[2];
    				Nready_in[2] = Sready_out[0];		
				end				
				
			end
	  	  end
   
  
    // ROUTER0
    Wdata_in[1]  = Edata_out[0];
    Wvalid_in[1] = Evalid_out[0];
    Eready_in[0] = Wready_out[1];
    Ndata_in[2]  = Sdata_out[0];
    Nvalid_in[2] = Svalid_out[0];
    Sready_in[0] = Nready_out[2];
    // ROUTER1
    Edata_in[0]  = Wdata_out[1];
    Evalid_in[0] = Wvalid_out[1];
    Wready_in[0] = Eready_out[0];
    Ndata_in[3]  = Sdata_out[1];
    Nvalid_in[3] = Svalid_out[1];
    Sready_in[1] = Nready_out[3];
    // ROUTER2
    Wdata_in[3]  = Edata_out[2];
    Wvalid_in[3] = Evalid_out[2];
    Eready_in[2] = Wready_out[3];
    Sdata_in[0]  = Ndata_out[2];
    Svalid_in[0] = Nvalid_out[2];
    Nready_in[2] = Sready_out[0];
    // ROUTER3
    Edata_in[2]  = Wdata_out[3];
    Evalid_in[2] = Wvalid_out[3];
    Wready_in[3] = Eready_out[2];
    Sdata_in[1]  = Ndata_out[3];
    Svalid_in[1] = Nvalid_out[3];
    Nready_in[3] = Sready_out[1];
  end
                  
  // Declaring the local variables
  reg [27 : 0]            data;               // 28 bits
  reg [2 : 0]             flit;
  reg                     parity = 1;
  reg [`DATA_WIDTH-1 : 0] tmp_data[`NODES-1 : 0];
  
  `include "tb_tasks_network.v"             // to include task predefined after declaring the signals
  
  // Specify the CYCLE parameter
  parameter CYCLE = 10;
  
  // Generating Clock of period 10ns
  initial begin
    clk = 0;
    forever 
      #(CYCLE/2) clk = ~clk;
  end
  
  // Start the simulation
  initial begin : SIM
    integer i;
    
    // Reset & Initialize
    // reset(.id, .Rxy_rst, .Cx_rst, .cur_addr_rst)
    // xpkt_gen(.id, .p_length, .d_addr, .s_addr, .p_id);
    reset('d0, 8'b00111100, 4'b1010, 4'b0000); //--NODE0
    reset('d1, 8'b00111100, 4'b1100, 4'b0001); //--NODE1
    reset('d2, 8'b00111100, 4'b0011, 4'b0010); //--NODE2
    reset('d3, 8'b00111100, 4'b0101, 4'b0011); //--NODE3
    Lpkt_gen('d3, 12'd5, 4'd0, 4'd3, 8'd5); // West
    Lpkt_gen('d2, 12'd6, 4'd0, 4'd2, 8'd6); // North
    fork
      Lpkt_gen('d0, 12'd4, 4'd3, 4'd0, 8'd4); // East
      Lpkt_gen('d2, 12'd7, 4'd0, 4'd2, 8'd7); // North
    join
    #(CYCLE * 25);
    $finish;
  end

endmodule